// cq_viola.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module cq_viola (
		input  wire        adc_MISO,      //      adc.MISO
		output wire        adc_MOSI,      //         .MOSI
		output wire        adc_SCLK,      //         .SCLK
		output wire        adc_SS_n,      //         .SS_n
		input  wire        clk_core_clk,  // clk_core.clk
		input  wire        clk_peri_clk,  // clk_peri.clk
		output wire        lcdc_rst_n,    //     lcdc.rst_n
		output wire        lcdc_cs_n,     //         .cs_n
		output wire        lcdc_rs,       //         .rs
		output wire        lcdc_wr_n,     //         .wr_n
		inout  wire [7:0]  lcdc_d,        //         .d
		output wire        led_export,    //      led.export
		output wire        mmc_nCS,       //      mmc.nCS
		output wire        mmc_SCK,       //         .SCK
		output wire        mmc_SDO,       //         .SDO
		input  wire        mmc_SDI,       //         .SDI
		input  wire        mmc_CD,        //         .CD
		input  wire        mmc_WP,        //         .WP
		input  wire        reset_reset_n, //    reset.reset_n
		output wire [11:0] sdr_addr,      //      sdr.addr
		output wire [1:0]  sdr_ba,        //         .ba
		output wire        sdr_cas_n,     //         .cas_n
		output wire        sdr_cke,       //         .cke
		output wire        sdr_cs_n,      //         .cs_n
		inout  wire [15:0] sdr_dq,        //         .dq
		output wire [1:0]  sdr_dqm,       //         .dqm
		output wire        sdr_ras_n,     //         .ras_n
		output wire        sdr_we_n,      //         .we_n
		output wire        sound_export   //    sound.export
	);

	wire  [31:0] nios2_s_custom_instruction_master_multi_dataa;                              // nios2_s:A_ci_multi_dataa -> nios2_s_custom_instruction_master_translator:ci_slave_multi_dataa
	wire         nios2_s_custom_instruction_master_multi_writerc;                            // nios2_s:A_ci_multi_writerc -> nios2_s_custom_instruction_master_translator:ci_slave_multi_writerc
	wire  [31:0] nios2_s_custom_instruction_master_multi_result;                             // nios2_s_custom_instruction_master_translator:ci_slave_multi_result -> nios2_s:A_ci_multi_result
	wire         nios2_s_custom_instruction_master_clk;                                      // nios2_s:A_ci_multi_clock -> nios2_s_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] nios2_s_custom_instruction_master_multi_datab;                              // nios2_s:A_ci_multi_datab -> nios2_s_custom_instruction_master_translator:ci_slave_multi_datab
	wire         nios2_s_custom_instruction_master_start;                                    // nios2_s:A_ci_multi_start -> nios2_s_custom_instruction_master_translator:ci_slave_multi_start
	wire   [4:0] nios2_s_custom_instruction_master_multi_b;                                  // nios2_s:A_ci_multi_b -> nios2_s_custom_instruction_master_translator:ci_slave_multi_b
	wire   [4:0] nios2_s_custom_instruction_master_multi_c;                                  // nios2_s:A_ci_multi_c -> nios2_s_custom_instruction_master_translator:ci_slave_multi_c
	wire         nios2_s_custom_instruction_master_reset_req;                                // nios2_s:A_ci_multi_reset_req -> nios2_s_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         nios2_s_custom_instruction_master_done;                                     // nios2_s_custom_instruction_master_translator:ci_slave_multi_done -> nios2_s:A_ci_multi_done
	wire   [4:0] nios2_s_custom_instruction_master_multi_a;                                  // nios2_s:A_ci_multi_a -> nios2_s_custom_instruction_master_translator:ci_slave_multi_a
	wire         nios2_s_custom_instruction_master_clk_en;                                   // nios2_s:A_ci_multi_clk_en -> nios2_s_custom_instruction_master_translator:ci_slave_multi_clken
	wire         nios2_s_custom_instruction_master_reset;                                    // nios2_s:A_ci_multi_reset -> nios2_s_custom_instruction_master_translator:ci_slave_multi_reset
	wire         nios2_s_custom_instruction_master_multi_readrb;                             // nios2_s:A_ci_multi_readrb -> nios2_s_custom_instruction_master_translator:ci_slave_multi_readrb
	wire         nios2_s_custom_instruction_master_multi_readra;                             // nios2_s:A_ci_multi_readra -> nios2_s_custom_instruction_master_translator:ci_slave_multi_readra
	wire   [7:0] nios2_s_custom_instruction_master_multi_n;                                  // nios2_s:A_ci_multi_n -> nios2_s_custom_instruction_master_translator:ci_slave_multi_n
	wire         nios2_s_custom_instruction_master_translator_multi_ci_master_readra;        // nios2_s_custom_instruction_master_translator:multi_ci_master_readra -> nios2_s_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] nios2_s_custom_instruction_master_translator_multi_ci_master_a;             // nios2_s_custom_instruction_master_translator:multi_ci_master_a -> nios2_s_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] nios2_s_custom_instruction_master_translator_multi_ci_master_b;             // nios2_s_custom_instruction_master_translator:multi_ci_master_b -> nios2_s_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         nios2_s_custom_instruction_master_translator_multi_ci_master_clk;           // nios2_s_custom_instruction_master_translator:multi_ci_master_clk -> nios2_s_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios2_s_custom_instruction_master_translator_multi_ci_master_readrb;        // nios2_s_custom_instruction_master_translator:multi_ci_master_readrb -> nios2_s_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] nios2_s_custom_instruction_master_translator_multi_ci_master_c;             // nios2_s_custom_instruction_master_translator:multi_ci_master_c -> nios2_s_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         nios2_s_custom_instruction_master_translator_multi_ci_master_start;         // nios2_s_custom_instruction_master_translator:multi_ci_master_start -> nios2_s_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         nios2_s_custom_instruction_master_translator_multi_ci_master_reset_req;     // nios2_s_custom_instruction_master_translator:multi_ci_master_reset_req -> nios2_s_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios2_s_custom_instruction_master_translator_multi_ci_master_done;          // nios2_s_custom_instruction_master_multi_xconnect:ci_slave_done -> nios2_s_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios2_s_custom_instruction_master_translator_multi_ci_master_n;             // nios2_s_custom_instruction_master_translator:multi_ci_master_n -> nios2_s_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] nios2_s_custom_instruction_master_translator_multi_ci_master_result;        // nios2_s_custom_instruction_master_multi_xconnect:ci_slave_result -> nios2_s_custom_instruction_master_translator:multi_ci_master_result
	wire         nios2_s_custom_instruction_master_translator_multi_ci_master_clk_en;        // nios2_s_custom_instruction_master_translator:multi_ci_master_clken -> nios2_s_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] nios2_s_custom_instruction_master_translator_multi_ci_master_datab;         // nios2_s_custom_instruction_master_translator:multi_ci_master_datab -> nios2_s_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] nios2_s_custom_instruction_master_translator_multi_ci_master_dataa;         // nios2_s_custom_instruction_master_translator:multi_ci_master_dataa -> nios2_s_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios2_s_custom_instruction_master_translator_multi_ci_master_reset;         // nios2_s_custom_instruction_master_translator:multi_ci_master_reset -> nios2_s_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         nios2_s_custom_instruction_master_translator_multi_ci_master_writerc;       // nios2_s_custom_instruction_master_translator:multi_ci_master_writerc -> nios2_s_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios2_s_custom_instruction_master_multi_xconnect_ci_master0_readra;         // nios2_s_custom_instruction_master_multi_xconnect:ci_master0_readra -> nios2_s_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_s_custom_instruction_master_multi_xconnect_ci_master0_a;              // nios2_s_custom_instruction_master_multi_xconnect:ci_master0_a -> nios2_s_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] nios2_s_custom_instruction_master_multi_xconnect_ci_master0_b;              // nios2_s_custom_instruction_master_multi_xconnect:ci_master0_b -> nios2_s_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         nios2_s_custom_instruction_master_multi_xconnect_ci_master0_readrb;         // nios2_s_custom_instruction_master_multi_xconnect:ci_master0_readrb -> nios2_s_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_s_custom_instruction_master_multi_xconnect_ci_master0_c;              // nios2_s_custom_instruction_master_multi_xconnect:ci_master0_c -> nios2_s_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios2_s_custom_instruction_master_multi_xconnect_ci_master0_clk;            // nios2_s_custom_instruction_master_multi_xconnect:ci_master0_clk -> nios2_s_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] nios2_s_custom_instruction_master_multi_xconnect_ci_master0_ipending;       // nios2_s_custom_instruction_master_multi_xconnect:ci_master0_ipending -> nios2_s_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios2_s_custom_instruction_master_multi_xconnect_ci_master0_start;          // nios2_s_custom_instruction_master_multi_xconnect:ci_master0_start -> nios2_s_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         nios2_s_custom_instruction_master_multi_xconnect_ci_master0_reset_req;      // nios2_s_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> nios2_s_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios2_s_custom_instruction_master_multi_xconnect_ci_master0_done;           // nios2_s_custom_instruction_master_multi_slave_translator0:ci_slave_done -> nios2_s_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] nios2_s_custom_instruction_master_multi_xconnect_ci_master0_n;              // nios2_s_custom_instruction_master_multi_xconnect:ci_master0_n -> nios2_s_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] nios2_s_custom_instruction_master_multi_xconnect_ci_master0_result;         // nios2_s_custom_instruction_master_multi_slave_translator0:ci_slave_result -> nios2_s_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         nios2_s_custom_instruction_master_multi_xconnect_ci_master0_estatus;        // nios2_s_custom_instruction_master_multi_xconnect:ci_master0_estatus -> nios2_s_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         nios2_s_custom_instruction_master_multi_xconnect_ci_master0_clk_en;         // nios2_s_custom_instruction_master_multi_xconnect:ci_master0_clken -> nios2_s_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] nios2_s_custom_instruction_master_multi_xconnect_ci_master0_datab;          // nios2_s_custom_instruction_master_multi_xconnect:ci_master0_datab -> nios2_s_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_s_custom_instruction_master_multi_xconnect_ci_master0_dataa;          // nios2_s_custom_instruction_master_multi_xconnect:ci_master0_dataa -> nios2_s_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios2_s_custom_instruction_master_multi_xconnect_ci_master0_reset;          // nios2_s_custom_instruction_master_multi_xconnect:ci_master0_reset -> nios2_s_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         nios2_s_custom_instruction_master_multi_xconnect_ci_master0_writerc;        // nios2_s_custom_instruction_master_multi_xconnect:ci_master0_writerc -> nios2_s_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_result; // pixelsimd:result -> nios2_s_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_clk;    // nios2_s_custom_instruction_master_multi_slave_translator0:ci_master_clk -> pixelsimd:clk
	wire         nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_clk_en; // nios2_s_custom_instruction_master_multi_slave_translator0:ci_master_clken -> pixelsimd:clk_en
	wire  [31:0] nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_datab;  // nios2_s_custom_instruction_master_multi_slave_translator0:ci_master_datab -> pixelsimd:datab
	wire  [31:0] nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_dataa;  // nios2_s_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> pixelsimd:dataa
	wire         nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_start;  // nios2_s_custom_instruction_master_multi_slave_translator0:ci_master_start -> pixelsimd:start
	wire         nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_reset;  // nios2_s_custom_instruction_master_multi_slave_translator0:ci_master_reset -> pixelsimd:reset
	wire         nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_done;   // pixelsimd:done -> nios2_s_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire   [2:0] nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_n;      // nios2_s_custom_instruction_master_multi_slave_translator0:ci_master_n -> pixelsimd:n
	wire  [31:0] nios2_s_data_master_readdata;                                               // mm_interconnect_0:nios2_s_data_master_readdata -> nios2_s:d_readdata
	wire         nios2_s_data_master_waitrequest;                                            // mm_interconnect_0:nios2_s_data_master_waitrequest -> nios2_s:d_waitrequest
	wire         nios2_s_data_master_debugaccess;                                            // nios2_s:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_s_data_master_debugaccess
	wire  [28:0] nios2_s_data_master_address;                                                // nios2_s:d_address -> mm_interconnect_0:nios2_s_data_master_address
	wire   [3:0] nios2_s_data_master_byteenable;                                             // nios2_s:d_byteenable -> mm_interconnect_0:nios2_s_data_master_byteenable
	wire         nios2_s_data_master_read;                                                   // nios2_s:d_read -> mm_interconnect_0:nios2_s_data_master_read
	wire         nios2_s_data_master_write;                                                  // nios2_s:d_write -> mm_interconnect_0:nios2_s_data_master_write
	wire  [31:0] nios2_s_data_master_writedata;                                              // nios2_s:d_writedata -> mm_interconnect_0:nios2_s_data_master_writedata
	wire  [31:0] nios2_s_instruction_master_readdata;                                        // mm_interconnect_0:nios2_s_instruction_master_readdata -> nios2_s:i_readdata
	wire         nios2_s_instruction_master_waitrequest;                                     // mm_interconnect_0:nios2_s_instruction_master_waitrequest -> nios2_s:i_waitrequest
	wire  [27:0] nios2_s_instruction_master_address;                                         // nios2_s:i_address -> mm_interconnect_0:nios2_s_instruction_master_address
	wire         nios2_s_instruction_master_read;                                            // nios2_s:i_read -> mm_interconnect_0:nios2_s_instruction_master_read
	wire         nios2_s_instruction_master_readdatavalid;                                   // mm_interconnect_0:nios2_s_instruction_master_readdatavalid -> nios2_s:i_readdatavalid
	wire   [3:0] nios2_s_instruction_master_burstcount;                                      // nios2_s:i_burstcount -> mm_interconnect_0:nios2_s_instruction_master_burstcount
	wire         lcdc_m1_waitrequest;                                                        // mm_interconnect_0:lcdc_m1_waitrequest -> lcdc:avm_m1_waitrequest
	wire  [15:0] lcdc_m1_readdata;                                                           // mm_interconnect_0:lcdc_m1_readdata -> lcdc:avm_m1_readdata
	wire  [30:0] lcdc_m1_address;                                                            // lcdc:avm_m1_address -> mm_interconnect_0:lcdc_m1_address
	wire         lcdc_m1_read;                                                               // lcdc:avm_m1_read -> mm_interconnect_0:lcdc_m1_read
	wire         lcdc_m1_readdatavalid;                                                      // mm_interconnect_0:lcdc_m1_readdatavalid -> lcdc:avm_m1_readdatavalid
	wire   [3:0] lcdc_m1_burstcount;                                                         // lcdc:avm_m1_burstcount -> mm_interconnect_0:lcdc_m1_burstcount
	wire  [31:0] mm_interconnect_0_nios2_s_debug_mem_slave_readdata;                         // nios2_s:debug_mem_slave_readdata -> mm_interconnect_0:nios2_s_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_s_debug_mem_slave_waitrequest;                      // nios2_s:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_s_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_s_debug_mem_slave_debugaccess;                      // mm_interconnect_0:nios2_s_debug_mem_slave_debugaccess -> nios2_s:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_s_debug_mem_slave_address;                          // mm_interconnect_0:nios2_s_debug_mem_slave_address -> nios2_s:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_s_debug_mem_slave_read;                             // mm_interconnect_0:nios2_s_debug_mem_slave_read -> nios2_s:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_s_debug_mem_slave_byteenable;                       // mm_interconnect_0:nios2_s_debug_mem_slave_byteenable -> nios2_s:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_s_debug_mem_slave_write;                            // mm_interconnect_0:nios2_s_debug_mem_slave_write -> nios2_s:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_s_debug_mem_slave_writedata;                        // mm_interconnect_0:nios2_s_debug_mem_slave_writedata -> nios2_s:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_mm_bridge_0_s0_readdata;                                  // mm_bridge_0:s0_readdata -> mm_interconnect_0:mm_bridge_0_s0_readdata
	wire         mm_interconnect_0_mm_bridge_0_s0_waitrequest;                               // mm_bridge_0:s0_waitrequest -> mm_interconnect_0:mm_bridge_0_s0_waitrequest
	wire         mm_interconnect_0_mm_bridge_0_s0_debugaccess;                               // mm_interconnect_0:mm_bridge_0_s0_debugaccess -> mm_bridge_0:s0_debugaccess
	wire  [15:0] mm_interconnect_0_mm_bridge_0_s0_address;                                   // mm_interconnect_0:mm_bridge_0_s0_address -> mm_bridge_0:s0_address
	wire         mm_interconnect_0_mm_bridge_0_s0_read;                                      // mm_interconnect_0:mm_bridge_0_s0_read -> mm_bridge_0:s0_read
	wire   [3:0] mm_interconnect_0_mm_bridge_0_s0_byteenable;                                // mm_interconnect_0:mm_bridge_0_s0_byteenable -> mm_bridge_0:s0_byteenable
	wire         mm_interconnect_0_mm_bridge_0_s0_readdatavalid;                             // mm_bridge_0:s0_readdatavalid -> mm_interconnect_0:mm_bridge_0_s0_readdatavalid
	wire         mm_interconnect_0_mm_bridge_0_s0_write;                                     // mm_interconnect_0:mm_bridge_0_s0_write -> mm_bridge_0:s0_write
	wire  [31:0] mm_interconnect_0_mm_bridge_0_s0_writedata;                                 // mm_interconnect_0:mm_bridge_0_s0_writedata -> mm_bridge_0:s0_writedata
	wire   [0:0] mm_interconnect_0_mm_bridge_0_s0_burstcount;                                // mm_interconnect_0:mm_bridge_0_s0_burstcount -> mm_bridge_0:s0_burstcount
	wire         mm_interconnect_0_sdram_s1_chipselect;                                      // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                        // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                     // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [21:0] mm_interconnect_0_sdram_s1_address;                                         // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                            // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                      // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                   // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                           // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                       // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_ipl_memory_s1_chipselect;                                 // mm_interconnect_0:ipl_memory_s1_chipselect -> ipl_memory:chipselect
	wire  [31:0] mm_interconnect_0_ipl_memory_s1_readdata;                                   // ipl_memory:readdata -> mm_interconnect_0:ipl_memory_s1_readdata
	wire  [10:0] mm_interconnect_0_ipl_memory_s1_address;                                    // mm_interconnect_0:ipl_memory_s1_address -> ipl_memory:address
	wire   [3:0] mm_interconnect_0_ipl_memory_s1_byteenable;                                 // mm_interconnect_0:ipl_memory_s1_byteenable -> ipl_memory:byteenable
	wire         mm_interconnect_0_ipl_memory_s1_write;                                      // mm_interconnect_0:ipl_memory_s1_write -> ipl_memory:write
	wire  [31:0] mm_interconnect_0_ipl_memory_s1_writedata;                                  // mm_interconnect_0:ipl_memory_s1_writedata -> ipl_memory:writedata
	wire         mm_interconnect_0_ipl_memory_s1_clken;                                      // mm_interconnect_0:ipl_memory_s1_clken -> ipl_memory:clken
	wire         mm_bridge_0_m0_waitrequest;                                                 // mm_interconnect_1:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	wire  [31:0] mm_bridge_0_m0_readdata;                                                    // mm_interconnect_1:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	wire         mm_bridge_0_m0_debugaccess;                                                 // mm_bridge_0:m0_debugaccess -> mm_interconnect_1:mm_bridge_0_m0_debugaccess
	wire  [15:0] mm_bridge_0_m0_address;                                                     // mm_bridge_0:m0_address -> mm_interconnect_1:mm_bridge_0_m0_address
	wire         mm_bridge_0_m0_read;                                                        // mm_bridge_0:m0_read -> mm_interconnect_1:mm_bridge_0_m0_read
	wire   [3:0] mm_bridge_0_m0_byteenable;                                                  // mm_bridge_0:m0_byteenable -> mm_interconnect_1:mm_bridge_0_m0_byteenable
	wire         mm_bridge_0_m0_readdatavalid;                                               // mm_interconnect_1:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	wire  [31:0] mm_bridge_0_m0_writedata;                                                   // mm_bridge_0:m0_writedata -> mm_interconnect_1:mm_bridge_0_m0_writedata
	wire         mm_bridge_0_m0_write;                                                       // mm_bridge_0:m0_write -> mm_interconnect_1:mm_bridge_0_m0_write
	wire   [0:0] mm_bridge_0_m0_burstcount;                                                  // mm_bridge_0:m0_burstcount -> mm_interconnect_1:mm_bridge_0_m0_burstcount
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;                   // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;                     // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest;                  // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;                      // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;                         // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;                        // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;                    // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;                             // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;                              // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire         mm_interconnect_1_systimer_s1_chipselect;                                   // mm_interconnect_1:systimer_s1_chipselect -> systimer:chipselect
	wire  [15:0] mm_interconnect_1_systimer_s1_readdata;                                     // systimer:readdata -> mm_interconnect_1:systimer_s1_readdata
	wire   [2:0] mm_interconnect_1_systimer_s1_address;                                      // mm_interconnect_1:systimer_s1_address -> systimer:address
	wire         mm_interconnect_1_systimer_s1_write;                                        // mm_interconnect_1:systimer_s1_write -> systimer:write_n
	wire  [15:0] mm_interconnect_1_systimer_s1_writedata;                                    // mm_interconnect_1:systimer_s1_writedata -> systimer:writedata
	wire         mm_interconnect_1_led_s1_chipselect;                                        // mm_interconnect_1:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_1_led_s1_readdata;                                          // led:readdata -> mm_interconnect_1:led_s1_readdata
	wire   [1:0] mm_interconnect_1_led_s1_address;                                           // mm_interconnect_1:led_s1_address -> led:address
	wire         mm_interconnect_1_led_s1_write;                                             // mm_interconnect_1:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_1_led_s1_writedata;                                         // mm_interconnect_1:led_s1_writedata -> led:writedata
	wire         mm_interconnect_1_mmcdma_s1_chipselect;                                     // mm_interconnect_1:mmcdma_s1_chipselect -> mmcdma:chipselect
	wire  [31:0] mm_interconnect_1_mmcdma_s1_readdata;                                       // mmcdma:readdata -> mm_interconnect_1:mmcdma_s1_readdata
	wire   [7:0] mm_interconnect_1_mmcdma_s1_address;                                        // mm_interconnect_1:mmcdma_s1_address -> mmcdma:address
	wire         mm_interconnect_1_mmcdma_s1_read;                                           // mm_interconnect_1:mmcdma_s1_read -> mmcdma:read
	wire         mm_interconnect_1_mmcdma_s1_write;                                          // mm_interconnect_1:mmcdma_s1_write -> mmcdma:write
	wire  [31:0] mm_interconnect_1_mmcdma_s1_writedata;                                      // mm_interconnect_1:mmcdma_s1_writedata -> mmcdma:writedata
	wire  [31:0] mm_interconnect_1_lcdc_s1_readdata;                                         // lcdc:avs_s1_readdata -> mm_interconnect_1:lcdc_s1_readdata
	wire   [1:0] mm_interconnect_1_lcdc_s1_address;                                          // mm_interconnect_1:lcdc_s1_address -> lcdc:avs_s1_address
	wire         mm_interconnect_1_lcdc_s1_read;                                             // mm_interconnect_1:lcdc_s1_read -> lcdc:avs_s1_read
	wire         mm_interconnect_1_lcdc_s1_write;                                            // mm_interconnect_1:lcdc_s1_write -> lcdc:avs_s1_write
	wire  [31:0] mm_interconnect_1_lcdc_s1_writedata;                                        // mm_interconnect_1:lcdc_s1_writedata -> lcdc:avs_s1_writedata
	wire   [7:0] mm_interconnect_1_sound_s1_readdata;                                        // sound:avs_s1_readdata -> mm_interconnect_1:sound_s1_readdata
	wire   [1:0] mm_interconnect_1_sound_s1_address;                                         // mm_interconnect_1:sound_s1_address -> sound:avs_s1_address
	wire         mm_interconnect_1_sound_s1_read;                                            // mm_interconnect_1:sound_s1_read -> sound:avs_s1_read
	wire         mm_interconnect_1_sound_s1_write;                                           // mm_interconnect_1:sound_s1_write -> sound:avs_s1_write
	wire   [7:0] mm_interconnect_1_sound_s1_writedata;                                       // mm_interconnect_1:sound_s1_writedata -> sound:avs_s1_writedata
	wire         mm_interconnect_1_touchpanel_spi_control_port_chipselect;                   // mm_interconnect_1:touchpanel_spi_control_port_chipselect -> touchpanel:spi_select
	wire  [15:0] mm_interconnect_1_touchpanel_spi_control_port_readdata;                     // touchpanel:data_to_cpu -> mm_interconnect_1:touchpanel_spi_control_port_readdata
	wire   [2:0] mm_interconnect_1_touchpanel_spi_control_port_address;                      // mm_interconnect_1:touchpanel_spi_control_port_address -> touchpanel:mem_addr
	wire         mm_interconnect_1_touchpanel_spi_control_port_read;                         // mm_interconnect_1:touchpanel_spi_control_port_read -> touchpanel:read_n
	wire         mm_interconnect_1_touchpanel_spi_control_port_write;                        // mm_interconnect_1:touchpanel_spi_control_port_write -> touchpanel:write_n
	wire  [15:0] mm_interconnect_1_touchpanel_spi_control_port_writedata;                    // mm_interconnect_1:touchpanel_spi_control_port_writedata -> touchpanel:data_from_cpu
	wire         irq_mapper_receiver1_irq;                                                   // lcdc:ins_s1_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_s_irq_irq;                                                            // irq_mapper:sender_irq -> nios2_s:irq
	wire         irq_mapper_receiver0_irq;                                                   // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                              // mmcdma:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver2_irq;                                                   // irq_synchronizer_001:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                                          // systimer:irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver3_irq;                                                   // irq_synchronizer_002:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                                          // jtag_uart:av_irq -> irq_synchronizer_002:receiver_irq
	wire         irq_mapper_receiver4_irq;                                                   // irq_synchronizer_003:sender_irq -> irq_mapper:receiver4_irq
	wire   [0:0] irq_synchronizer_003_receiver_irq;                                          // touchpanel:irq -> irq_synchronizer_003:receiver_irq
	wire         irq_mapper_receiver5_irq;                                                   // irq_synchronizer_004:sender_irq -> irq_mapper:receiver5_irq
	wire   [0:0] irq_synchronizer_004_receiver_irq;                                          // sound:avs_s1_irq -> irq_synchronizer_004:receiver_irq
	wire         rst_controller_reset_out_reset;                                             // rst_controller:reset_out -> [ipl_memory:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, lcdc:csi_reset, mm_interconnect_0:nios2_s_reset_reset_bridge_in_reset_reset, mm_interconnect_1:lcdc_clock_reset_reset_bridge_in_reset_reset, nios2_s:reset_n, rst_translator:in_reset, sdram:reset_n]
	wire         rst_controller_reset_out_reset_req;                                         // rst_controller:reset_req -> [ipl_memory:reset_req, nios2_s:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                         // rst_controller_001:reset_out -> [irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, irq_synchronizer_004:receiver_reset, jtag_uart:rst_n, led:reset_n, mm_bridge_0:reset, mm_interconnect_0:mm_bridge_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:mm_bridge_0_reset_reset_bridge_in_reset_reset, mmcdma:reset, sound:csi_global_reset, sysid:reset_n, systimer:reset_n, touchpanel:reset_n]

	cq_viola_ipl_memory ipl_memory (
		.clk        (clk_core_clk),                               //   clk1.clk
		.address    (mm_interconnect_0_ipl_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ipl_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ipl_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ipl_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ipl_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ipl_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ipl_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)          //       .reset_req
	);

	cq_viola_jtag_uart jtag_uart (
		.clk            (clk_peri_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_002_receiver_irq)                          //               irq.irq
	);

	lcdc_component lcdc (
		.csi_clk              (clk_core_clk),                        //            clock.clk
		.csi_reset            (rst_controller_reset_out_reset),      //      clock_reset.reset
		.avs_s1_address       (mm_interconnect_1_lcdc_s1_address),   //               s1.address
		.avs_s1_read          (mm_interconnect_1_lcdc_s1_read),      //                 .read
		.avs_s1_readdata      (mm_interconnect_1_lcdc_s1_readdata),  //                 .readdata
		.avs_s1_write         (mm_interconnect_1_lcdc_s1_write),     //                 .write
		.avs_s1_writedata     (mm_interconnect_1_lcdc_s1_writedata), //                 .writedata
		.avm_m1_address       (lcdc_m1_address),                     //               m1.address
		.avm_m1_waitrequest   (lcdc_m1_waitrequest),                 //                 .waitrequest
		.avm_m1_burstcount    (lcdc_m1_burstcount),                  //                 .burstcount
		.avm_m1_read          (lcdc_m1_read),                        //                 .read
		.avm_m1_readdata      (lcdc_m1_readdata),                    //                 .readdata
		.avm_m1_readdatavalid (lcdc_m1_readdatavalid),               //                 .readdatavalid
		.coe_lcd_rst_n        (lcdc_rst_n),                          //    conduit_end_0.export
		.coe_lcd_cs_n         (lcdc_cs_n),                           //                 .export
		.coe_lcd_rs           (lcdc_rs),                             //                 .export
		.coe_lcd_wr_n         (lcdc_wr_n),                           //                 .export
		.coe_lcd_d            (lcdc_d),                              //                 .export
		.ins_s1_irq           (irq_mapper_receiver1_irq)             // interrupt_sender.irq
	);

	cq_viola_led led (
		.clk        (clk_peri_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                           // external_connection.export
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (16),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_0 (
		.clk              (clk_peri_clk),                                   //   clk.clk
		.reset            (rst_controller_001_reset_out_reset),             // reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_bridge_0_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_bridge_0_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_bridge_0_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_bridge_0_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_mm_bridge_0_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_mm_bridge_0_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_mm_bridge_0_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_mm_bridge_0_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_mm_bridge_0_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_bridge_0_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_0_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_0_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_0_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_0_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_0_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_0_m0_address),                         //      .address
		.m0_write         (mm_bridge_0_m0_write),                           //      .write
		.m0_read          (mm_bridge_0_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_0_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_0_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                               // (terminated)
		.m0_response      (2'b00)                                           // (terminated)
	);

	avalonif_mmcdma #(
		.SYSTEMCLOCKINFO (40000000)
	) mmcdma (
		.clk        (clk_peri_clk),                           //       clock_reset.clk
		.reset      (rst_controller_001_reset_out_reset),     // clock_reset_reset.reset
		.chipselect (mm_interconnect_1_mmcdma_s1_chipselect), //                s1.chipselect
		.address    (mm_interconnect_1_mmcdma_s1_address),    //                  .address
		.read       (mm_interconnect_1_mmcdma_s1_read),       //                  .read
		.readdata   (mm_interconnect_1_mmcdma_s1_readdata),   //                  .readdata
		.write      (mm_interconnect_1_mmcdma_s1_write),      //                  .write
		.writedata  (mm_interconnect_1_mmcdma_s1_writedata),  //                  .writedata
		.MMC_nCS    (mmc_nCS),                                //       conduit_end.export
		.MMC_SCK    (mmc_SCK),                                //                  .export
		.MMC_SDO    (mmc_SDO),                                //                  .export
		.MMC_SDI    (mmc_SDI),                                //                  .export
		.MMC_CD     (mmc_CD),                                 //                  .export
		.MMC_WP     (mmc_WP),                                 //                  .export
		.irq        (irq_synchronizer_receiver_irq)           //  interrupt_sender.irq
	);

	cq_viola_nios2_s nios2_s (
		.clk                                 (clk_core_clk),                                          //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                       //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                           (nios2_s_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_s_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_s_data_master_read),                              //                          .read
		.d_readdata                          (nios2_s_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_s_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_s_data_master_write),                             //                          .write
		.d_writedata                         (nios2_s_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_s_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_s_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_s_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_s_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_s_instruction_master_waitrequest),                //                          .waitrequest
		.i_burstcount                        (nios2_s_instruction_master_burstcount),                 //                          .burstcount
		.i_readdatavalid                     (nios2_s_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_s_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                      //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_s_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_s_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_s_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_s_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_s_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_s_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_s_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_s_debug_mem_slave_writedata),   //                          .writedata
		.A_ci_multi_done                     (nios2_s_custom_instruction_master_done),                // custom_instruction_master.done
		.A_ci_multi_result                   (nios2_s_custom_instruction_master_multi_result),        //                          .multi_result
		.A_ci_multi_a                        (nios2_s_custom_instruction_master_multi_a),             //                          .multi_a
		.A_ci_multi_b                        (nios2_s_custom_instruction_master_multi_b),             //                          .multi_b
		.A_ci_multi_c                        (nios2_s_custom_instruction_master_multi_c),             //                          .multi_c
		.A_ci_multi_clk_en                   (nios2_s_custom_instruction_master_clk_en),              //                          .clk_en
		.A_ci_multi_clock                    (nios2_s_custom_instruction_master_clk),                 //                          .clk
		.A_ci_multi_reset                    (nios2_s_custom_instruction_master_reset),               //                          .reset
		.A_ci_multi_reset_req                (nios2_s_custom_instruction_master_reset_req),           //                          .reset_req
		.A_ci_multi_dataa                    (nios2_s_custom_instruction_master_multi_dataa),         //                          .multi_dataa
		.A_ci_multi_datab                    (nios2_s_custom_instruction_master_multi_datab),         //                          .multi_datab
		.A_ci_multi_n                        (nios2_s_custom_instruction_master_multi_n),             //                          .multi_n
		.A_ci_multi_readra                   (nios2_s_custom_instruction_master_multi_readra),        //                          .multi_readra
		.A_ci_multi_readrb                   (nios2_s_custom_instruction_master_multi_readrb),        //                          .multi_readrb
		.A_ci_multi_start                    (nios2_s_custom_instruction_master_start),               //                          .start
		.A_ci_multi_writerc                  (nios2_s_custom_instruction_master_multi_writerc)        //                          .multi_writerc
	);

	pixelsimd pixelsimd (
		.dataa  (nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // nios_custom_instruction_slave_0.dataa
		.datab  (nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //                                .datab
		.result (nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_result), //                                .result
		.clk    (nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //                                .clk
		.clk_en (nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //                                .clk_en
		.reset  (nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //                                .reset
		.start  (nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_start),  //                                .start
		.done   (nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_done),   //                                .done
		.n      (nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_n)       //                                .n
	);

	cq_viola_sdram sdram (
		.clk            (clk_core_clk),                             //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdr_addr),                                 //  wire.export
		.zs_ba          (sdr_ba),                                   //      .export
		.zs_cas_n       (sdr_cas_n),                                //      .export
		.zs_cke         (sdr_cke),                                  //      .export
		.zs_cs_n        (sdr_cs_n),                                 //      .export
		.zs_dq          (sdr_dq),                                   //      .export
		.zs_dqm         (sdr_dqm),                                  //      .export
		.zs_ras_n       (sdr_ras_n),                                //      .export
		.zs_we_n        (sdr_we_n)                                  //      .export
	);

	avalonif_sound sound (
		.csi_global_clk   (clk_peri_clk),                         //       global.clk
		.csi_global_reset (rst_controller_001_reset_out_reset),   // global_reset.reset
		.avs_s1_address   (mm_interconnect_1_sound_s1_address),   //           s1.address
		.avs_s1_read      (mm_interconnect_1_sound_s1_read),      //             .read
		.avs_s1_readdata  (mm_interconnect_1_sound_s1_readdata),  //             .readdata
		.avs_s1_write     (mm_interconnect_1_sound_s1_write),     //             .write
		.avs_s1_writedata (mm_interconnect_1_sound_s1_writedata), //             .writedata
		.avs_s1_irq       (irq_synchronizer_004_receiver_irq),    //       irq_s1.irq
		.dac_out          (sound_export)                          //  conduit_end.export
	);

	cq_viola_sysid sysid (
		.clock    (clk_peri_clk),                                   //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	cq_viola_systimer systimer (
		.clk        (clk_peri_clk),                             //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.address    (mm_interconnect_1_systimer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_systimer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_systimer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_systimer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_systimer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_001_receiver_irq)         //   irq.irq
	);

	cq_viola_touchpanel touchpanel (
		.clk           (clk_peri_clk),                                             //              clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                      //            reset.reset_n
		.data_from_cpu (mm_interconnect_1_touchpanel_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_1_touchpanel_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_1_touchpanel_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_1_touchpanel_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_1_touchpanel_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_1_touchpanel_spi_control_port_write),     //                 .write_n
		.irq           (irq_synchronizer_003_receiver_irq),                        //              irq.irq
		.MISO          (adc_MISO),                                                 //         external.export
		.MOSI          (adc_MOSI),                                                 //                 .export
		.SCLK          (adc_SCLK),                                                 //                 .export
		.SS_n          (adc_SS_n)                                                  //                 .export
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) nios2_s_custom_instruction_master_translator (
		.ci_slave_result           (),                                                                       //        ci_slave.result
		.ci_slave_multi_clk        (nios2_s_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios2_s_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios2_s_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios2_s_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios2_s_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios2_s_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (nios2_s_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (nios2_s_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (nios2_s_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (nios2_s_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (nios2_s_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (nios2_s_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (nios2_s_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (nios2_s_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (nios2_s_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (nios2_s_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_result     (),                                                                       //  comb_ci_master.result
		.multi_ci_master_clk       (nios2_s_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios2_s_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios2_s_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios2_s_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios2_s_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios2_s_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios2_s_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios2_s_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios2_s_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios2_s_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios2_s_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios2_s_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios2_s_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios2_s_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios2_s_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios2_s_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_dataa            (32'b00000000000000000000000000000000),                                   //     (terminated)
		.ci_slave_datab            (32'b00000000000000000000000000000000),                                   //     (terminated)
		.ci_slave_n                (8'b00000000),                                                            //     (terminated)
		.ci_slave_readra           (1'b0),                                                                   //     (terminated)
		.ci_slave_readrb           (1'b0),                                                                   //     (terminated)
		.ci_slave_writerc          (1'b0),                                                                   //     (terminated)
		.ci_slave_a                (5'b00000),                                                               //     (terminated)
		.ci_slave_b                (5'b00000),                                                               //     (terminated)
		.ci_slave_c                (5'b00000),                                                               //     (terminated)
		.ci_slave_ipending         (32'b00000000000000000000000000000000),                                   //     (terminated)
		.ci_slave_estatus          (1'b0),                                                                   //     (terminated)
		.comb_ci_master_dataa      (),                                                                       //     (terminated)
		.comb_ci_master_datab      (),                                                                       //     (terminated)
		.comb_ci_master_n          (),                                                                       //     (terminated)
		.comb_ci_master_readra     (),                                                                       //     (terminated)
		.comb_ci_master_readrb     (),                                                                       //     (terminated)
		.comb_ci_master_writerc    (),                                                                       //     (terminated)
		.comb_ci_master_a          (),                                                                       //     (terminated)
		.comb_ci_master_b          (),                                                                       //     (terminated)
		.comb_ci_master_c          (),                                                                       //     (terminated)
		.comb_ci_master_ipending   (),                                                                       //     (terminated)
		.comb_ci_master_estatus    ()                                                                        //     (terminated)
	);

	cq_viola_nios2_s_custom_instruction_master_multi_xconnect nios2_s_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios2_s_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios2_s_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios2_s_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios2_s_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios2_s_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios2_s_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios2_s_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios2_s_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios2_s_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios2_s_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                       //           .ipending
		.ci_slave_estatus     (),                                                                       //           .estatus
		.ci_slave_clk         (nios2_s_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios2_s_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios2_s_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios2_s_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios2_s_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios2_s_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios2_s_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (nios2_s_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_n),      //          .n
		.ci_master_clk       (nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (nios2_s_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_readra    (),                                                                           // (terminated)
		.ci_master_readrb    (),                                                                           // (terminated)
		.ci_master_writerc   (),                                                                           // (terminated)
		.ci_master_a         (),                                                                           // (terminated)
		.ci_master_b         (),                                                                           // (terminated)
		.ci_master_c         (),                                                                           // (terminated)
		.ci_master_ipending  (),                                                                           // (terminated)
		.ci_master_estatus   (),                                                                           // (terminated)
		.ci_master_reset_req ()                                                                            // (terminated)
	);

	cq_viola_mm_interconnect_0 mm_interconnect_0 (
		.clk_core_clk_clk                              (clk_core_clk),                                          //                            clk_core_clk.clk
		.clk_peri_clk_clk                              (clk_peri_clk),                                          //                            clk_peri_clk.clk
		.mm_bridge_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                    // mm_bridge_0_reset_reset_bridge_in_reset.reset
		.nios2_s_reset_reset_bridge_in_reset_reset     (rst_controller_reset_out_reset),                        //     nios2_s_reset_reset_bridge_in_reset.reset
		.lcdc_m1_address                               (lcdc_m1_address),                                       //                                 lcdc_m1.address
		.lcdc_m1_waitrequest                           (lcdc_m1_waitrequest),                                   //                                        .waitrequest
		.lcdc_m1_burstcount                            (lcdc_m1_burstcount),                                    //                                        .burstcount
		.lcdc_m1_read                                  (lcdc_m1_read),                                          //                                        .read
		.lcdc_m1_readdata                              (lcdc_m1_readdata),                                      //                                        .readdata
		.lcdc_m1_readdatavalid                         (lcdc_m1_readdatavalid),                                 //                                        .readdatavalid
		.nios2_s_data_master_address                   (nios2_s_data_master_address),                           //                     nios2_s_data_master.address
		.nios2_s_data_master_waitrequest               (nios2_s_data_master_waitrequest),                       //                                        .waitrequest
		.nios2_s_data_master_byteenable                (nios2_s_data_master_byteenable),                        //                                        .byteenable
		.nios2_s_data_master_read                      (nios2_s_data_master_read),                              //                                        .read
		.nios2_s_data_master_readdata                  (nios2_s_data_master_readdata),                          //                                        .readdata
		.nios2_s_data_master_write                     (nios2_s_data_master_write),                             //                                        .write
		.nios2_s_data_master_writedata                 (nios2_s_data_master_writedata),                         //                                        .writedata
		.nios2_s_data_master_debugaccess               (nios2_s_data_master_debugaccess),                       //                                        .debugaccess
		.nios2_s_instruction_master_address            (nios2_s_instruction_master_address),                    //              nios2_s_instruction_master.address
		.nios2_s_instruction_master_waitrequest        (nios2_s_instruction_master_waitrequest),                //                                        .waitrequest
		.nios2_s_instruction_master_burstcount         (nios2_s_instruction_master_burstcount),                 //                                        .burstcount
		.nios2_s_instruction_master_read               (nios2_s_instruction_master_read),                       //                                        .read
		.nios2_s_instruction_master_readdata           (nios2_s_instruction_master_readdata),                   //                                        .readdata
		.nios2_s_instruction_master_readdatavalid      (nios2_s_instruction_master_readdatavalid),              //                                        .readdatavalid
		.ipl_memory_s1_address                         (mm_interconnect_0_ipl_memory_s1_address),               //                           ipl_memory_s1.address
		.ipl_memory_s1_write                           (mm_interconnect_0_ipl_memory_s1_write),                 //                                        .write
		.ipl_memory_s1_readdata                        (mm_interconnect_0_ipl_memory_s1_readdata),              //                                        .readdata
		.ipl_memory_s1_writedata                       (mm_interconnect_0_ipl_memory_s1_writedata),             //                                        .writedata
		.ipl_memory_s1_byteenable                      (mm_interconnect_0_ipl_memory_s1_byteenable),            //                                        .byteenable
		.ipl_memory_s1_chipselect                      (mm_interconnect_0_ipl_memory_s1_chipselect),            //                                        .chipselect
		.ipl_memory_s1_clken                           (mm_interconnect_0_ipl_memory_s1_clken),                 //                                        .clken
		.mm_bridge_0_s0_address                        (mm_interconnect_0_mm_bridge_0_s0_address),              //                          mm_bridge_0_s0.address
		.mm_bridge_0_s0_write                          (mm_interconnect_0_mm_bridge_0_s0_write),                //                                        .write
		.mm_bridge_0_s0_read                           (mm_interconnect_0_mm_bridge_0_s0_read),                 //                                        .read
		.mm_bridge_0_s0_readdata                       (mm_interconnect_0_mm_bridge_0_s0_readdata),             //                                        .readdata
		.mm_bridge_0_s0_writedata                      (mm_interconnect_0_mm_bridge_0_s0_writedata),            //                                        .writedata
		.mm_bridge_0_s0_burstcount                     (mm_interconnect_0_mm_bridge_0_s0_burstcount),           //                                        .burstcount
		.mm_bridge_0_s0_byteenable                     (mm_interconnect_0_mm_bridge_0_s0_byteenable),           //                                        .byteenable
		.mm_bridge_0_s0_readdatavalid                  (mm_interconnect_0_mm_bridge_0_s0_readdatavalid),        //                                        .readdatavalid
		.mm_bridge_0_s0_waitrequest                    (mm_interconnect_0_mm_bridge_0_s0_waitrequest),          //                                        .waitrequest
		.mm_bridge_0_s0_debugaccess                    (mm_interconnect_0_mm_bridge_0_s0_debugaccess),          //                                        .debugaccess
		.nios2_s_debug_mem_slave_address               (mm_interconnect_0_nios2_s_debug_mem_slave_address),     //                 nios2_s_debug_mem_slave.address
		.nios2_s_debug_mem_slave_write                 (mm_interconnect_0_nios2_s_debug_mem_slave_write),       //                                        .write
		.nios2_s_debug_mem_slave_read                  (mm_interconnect_0_nios2_s_debug_mem_slave_read),        //                                        .read
		.nios2_s_debug_mem_slave_readdata              (mm_interconnect_0_nios2_s_debug_mem_slave_readdata),    //                                        .readdata
		.nios2_s_debug_mem_slave_writedata             (mm_interconnect_0_nios2_s_debug_mem_slave_writedata),   //                                        .writedata
		.nios2_s_debug_mem_slave_byteenable            (mm_interconnect_0_nios2_s_debug_mem_slave_byteenable),  //                                        .byteenable
		.nios2_s_debug_mem_slave_waitrequest           (mm_interconnect_0_nios2_s_debug_mem_slave_waitrequest), //                                        .waitrequest
		.nios2_s_debug_mem_slave_debugaccess           (mm_interconnect_0_nios2_s_debug_mem_slave_debugaccess), //                                        .debugaccess
		.sdram_s1_address                              (mm_interconnect_0_sdram_s1_address),                    //                                sdram_s1.address
		.sdram_s1_write                                (mm_interconnect_0_sdram_s1_write),                      //                                        .write
		.sdram_s1_read                                 (mm_interconnect_0_sdram_s1_read),                       //                                        .read
		.sdram_s1_readdata                             (mm_interconnect_0_sdram_s1_readdata),                   //                                        .readdata
		.sdram_s1_writedata                            (mm_interconnect_0_sdram_s1_writedata),                  //                                        .writedata
		.sdram_s1_byteenable                           (mm_interconnect_0_sdram_s1_byteenable),                 //                                        .byteenable
		.sdram_s1_readdatavalid                        (mm_interconnect_0_sdram_s1_readdatavalid),              //                                        .readdatavalid
		.sdram_s1_waitrequest                          (mm_interconnect_0_sdram_s1_waitrequest),                //                                        .waitrequest
		.sdram_s1_chipselect                           (mm_interconnect_0_sdram_s1_chipselect)                  //                                        .chipselect
	);

	cq_viola_mm_interconnect_1 mm_interconnect_1 (
		.clk_core_clk_clk                              (clk_core_clk),                                              //                            clk_core_clk.clk
		.clk_peri_clk_clk                              (clk_peri_clk),                                              //                            clk_peri_clk.clk
		.lcdc_clock_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                            //  lcdc_clock_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                        // mm_bridge_0_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_m0_address                        (mm_bridge_0_m0_address),                                    //                          mm_bridge_0_m0.address
		.mm_bridge_0_m0_waitrequest                    (mm_bridge_0_m0_waitrequest),                                //                                        .waitrequest
		.mm_bridge_0_m0_burstcount                     (mm_bridge_0_m0_burstcount),                                 //                                        .burstcount
		.mm_bridge_0_m0_byteenable                     (mm_bridge_0_m0_byteenable),                                 //                                        .byteenable
		.mm_bridge_0_m0_read                           (mm_bridge_0_m0_read),                                       //                                        .read
		.mm_bridge_0_m0_readdata                       (mm_bridge_0_m0_readdata),                                   //                                        .readdata
		.mm_bridge_0_m0_readdatavalid                  (mm_bridge_0_m0_readdatavalid),                              //                                        .readdatavalid
		.mm_bridge_0_m0_write                          (mm_bridge_0_m0_write),                                      //                                        .write
		.mm_bridge_0_m0_writedata                      (mm_bridge_0_m0_writedata),                                  //                                        .writedata
		.mm_bridge_0_m0_debugaccess                    (mm_bridge_0_m0_debugaccess),                                //                                        .debugaccess
		.jtag_uart_avalon_jtag_slave_address           (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //             jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write             (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),       //                                        .write
		.jtag_uart_avalon_jtag_slave_read              (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),        //                                        .read
		.jtag_uart_avalon_jtag_slave_readdata          (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                                        .readdata
		.jtag_uart_avalon_jtag_slave_writedata         (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                                        .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest       (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                                        .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect        (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  //                                        .chipselect
		.lcdc_s1_address                               (mm_interconnect_1_lcdc_s1_address),                         //                                 lcdc_s1.address
		.lcdc_s1_write                                 (mm_interconnect_1_lcdc_s1_write),                           //                                        .write
		.lcdc_s1_read                                  (mm_interconnect_1_lcdc_s1_read),                            //                                        .read
		.lcdc_s1_readdata                              (mm_interconnect_1_lcdc_s1_readdata),                        //                                        .readdata
		.lcdc_s1_writedata                             (mm_interconnect_1_lcdc_s1_writedata),                       //                                        .writedata
		.led_s1_address                                (mm_interconnect_1_led_s1_address),                          //                                  led_s1.address
		.led_s1_write                                  (mm_interconnect_1_led_s1_write),                            //                                        .write
		.led_s1_readdata                               (mm_interconnect_1_led_s1_readdata),                         //                                        .readdata
		.led_s1_writedata                              (mm_interconnect_1_led_s1_writedata),                        //                                        .writedata
		.led_s1_chipselect                             (mm_interconnect_1_led_s1_chipselect),                       //                                        .chipselect
		.mmcdma_s1_address                             (mm_interconnect_1_mmcdma_s1_address),                       //                               mmcdma_s1.address
		.mmcdma_s1_write                               (mm_interconnect_1_mmcdma_s1_write),                         //                                        .write
		.mmcdma_s1_read                                (mm_interconnect_1_mmcdma_s1_read),                          //                                        .read
		.mmcdma_s1_readdata                            (mm_interconnect_1_mmcdma_s1_readdata),                      //                                        .readdata
		.mmcdma_s1_writedata                           (mm_interconnect_1_mmcdma_s1_writedata),                     //                                        .writedata
		.mmcdma_s1_chipselect                          (mm_interconnect_1_mmcdma_s1_chipselect),                    //                                        .chipselect
		.sound_s1_address                              (mm_interconnect_1_sound_s1_address),                        //                                sound_s1.address
		.sound_s1_write                                (mm_interconnect_1_sound_s1_write),                          //                                        .write
		.sound_s1_read                                 (mm_interconnect_1_sound_s1_read),                           //                                        .read
		.sound_s1_readdata                             (mm_interconnect_1_sound_s1_readdata),                       //                                        .readdata
		.sound_s1_writedata                            (mm_interconnect_1_sound_s1_writedata),                      //                                        .writedata
		.sysid_control_slave_address                   (mm_interconnect_1_sysid_control_slave_address),             //                     sysid_control_slave.address
		.sysid_control_slave_readdata                  (mm_interconnect_1_sysid_control_slave_readdata),            //                                        .readdata
		.systimer_s1_address                           (mm_interconnect_1_systimer_s1_address),                     //                             systimer_s1.address
		.systimer_s1_write                             (mm_interconnect_1_systimer_s1_write),                       //                                        .write
		.systimer_s1_readdata                          (mm_interconnect_1_systimer_s1_readdata),                    //                                        .readdata
		.systimer_s1_writedata                         (mm_interconnect_1_systimer_s1_writedata),                   //                                        .writedata
		.systimer_s1_chipselect                        (mm_interconnect_1_systimer_s1_chipselect),                  //                                        .chipselect
		.touchpanel_spi_control_port_address           (mm_interconnect_1_touchpanel_spi_control_port_address),     //             touchpanel_spi_control_port.address
		.touchpanel_spi_control_port_write             (mm_interconnect_1_touchpanel_spi_control_port_write),       //                                        .write
		.touchpanel_spi_control_port_read              (mm_interconnect_1_touchpanel_spi_control_port_read),        //                                        .read
		.touchpanel_spi_control_port_readdata          (mm_interconnect_1_touchpanel_spi_control_port_readdata),    //                                        .readdata
		.touchpanel_spi_control_port_writedata         (mm_interconnect_1_touchpanel_spi_control_port_writedata),   //                                        .writedata
		.touchpanel_spi_control_port_chipselect        (mm_interconnect_1_touchpanel_spi_control_port_chipselect)   //                                        .chipselect
	);

	cq_viola_irq_mapper irq_mapper (
		.clk           (clk_core_clk),                   //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.sender_irq    (nios2_s_irq_irq)                 //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_peri_clk),                       //       receiver_clk.clk
		.sender_clk     (clk_core_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk_peri_clk),                       //       receiver_clk.clk
		.sender_clk     (clk_core_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (clk_peri_clk),                       //       receiver_clk.clk
		.sender_clk     (clk_core_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (clk_peri_clk),                       //       receiver_clk.clk
		.sender_clk     (clk_core_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_004 (
		.receiver_clk   (clk_peri_clk),                       //       receiver_clk.clk
		.sender_clk     (clk_core_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_004_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver5_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_core_clk),                       //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_peri_clk),                       //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
